VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS	1000 ;
END UNITS

MANUFACTURINGGRID	0.005 ;

SITE core
  SIZE 0.20 BY 2.00 ;
  CLASS CORE ;
END core

LAYER metal1
  TYPE			ROUTING ;
  DIRECTION		HORIZONTAL ;
  PITCH			0.200 ;
  OFFSET		0.000 ;
  WIDTH			0.100 ;
END metal1

LAYER metal2
  TYPE			ROUTING ;
  DIRECTION		VERTICAL ;
  PITCH			0.200 ;
  OFFSET		0.100 ;
  WIDTH			0.1 ;
END metal2

LAYER metal3
  TYPE			ROUTING ;
  DIRECTION		HORIZONTAL ;
  PITCH			0.200 ;
  OFFSET		0.000 ;
  WIDTH			0.1 ;
END metal3

MACRO DFF_X1
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.6 BY 2.0 ;

  SITE  core ;
  PIN Q DIRECTION OUTPUT ;
    PORT
			LAYER metal2 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END Q 
  PIN CK DIRECTION INPUT ;
    PORT
			LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END CK
  PIN D DIRECTION INPUT ;
    PORT
			LAYER metal1 ;
      RECT 1.05 0.500 1.15 1.500 ;
    END
  END D
END DFF_X1 

MACRO INV_X1
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 0.8 BY 2.0 ;

  SITE  core ;
  PIN ZN DIRECTION OUTPUT ;
    PORT
			LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END ZN
  PIN A DIRECTION INPUT ;
    PORT
			LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END A
END INV_X1

MACRO INV_X8
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 6.4 BY 2.0 ;

  SITE  core ;
  PIN ZN DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END ZN
  PIN A DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
      RECT 3.25 0.500 3.35 1.500 ;
    END
  END A
END INV_X8

MACRO NAND2_X1
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;

  SITE  core ;
  PIN ZN DIRECTION OUTPUT ;
    PORT
			LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END ZN 
  PIN A1 DIRECTION INPUT ;
    PORT
			LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END A1
  PIN A2 DIRECTION INPUT ;
    PORT
			LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END A2
END NAND2_X1

MACRO NOR2_X1
  CLASS CORE ;
  ORIGIN 0 0  ;
  SIZE 1.2 BY 2.0 ;

  SITE  core ;
  PIN ZN DIRECTION OUTPUT ;
    PORT
			LAYER metal1 ;
      RECT 0.05 0.500 0.15 1.500 ;
    END
  END ZN
  PIN A1 DIRECTION INPUT ;
    PORT
			LAYER metal1 ;
      RECT 0.45 0.500 0.55 1.500 ;
    END
  END A1
  PIN A2 DIRECTION INPUT ;
    PORT
			LAYER metal1 ;
      RECT 0.85 0.500 0.95 1.500 ;
    END
  END A2
END NOR2_X1

END LIBRARY
